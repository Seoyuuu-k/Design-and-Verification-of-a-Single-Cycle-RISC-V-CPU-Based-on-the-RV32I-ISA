// `timescale 1ns / 1ps

// //rom
module instr_mem (
    input  logic [31:0] instr_rAddr,
    output logic [31:0] instr_code
);
    logic [31:0] rom [0:128];

initial begin
    // $readmemh("code2.txt",rom);
     $readmemh("code_mem.mem",rom);
end
// //---------------------------------------------------------------------------------------------------------------//
// //--------------------------------------------for_Rtype----------------------------------------------------------//
// //---------------------------------------------------------------------------------------------------------------//

//       initial begin
//     // add x11, x3, x4 -> x11 = 3 + 4 = 7
//     rom[0] = 32'h004185B3; 
//     // sub x2, x2, x1    -> x2 = 2 - 1 = 1
//     rom[1]  = 32'h40110133;
//     // and x4, x5, x4    -> 5 & 4 = 4
//     rom[2]  = 32'h0042F233; 
//     // or x3, x5, x4     -> 5 | 4 = 5
//     rom[3]  = 32'h0042E1B3; 
//     // xor x7, x5, x4    -> 5 ^ 4 = 1
//     rom[4]  = 32'h0042C3B3; 
//     // sll x4, x4, x7    -> 4 << 1 = 8
//     rom[5]  = 32'h00721233; 
//     // srl x3, x3, x7    -> 5 >> 1 = 2
//     rom[6]  = 32'h0071D1B3; 
//     // sra x9, x9, x7    -> (sign extend) >> 1
//     // sra (sign) msb 1 // x9== 32'b1100000....;
//     rom[7]  = 32'h4074D4B3; 
//     // sra x8, x8, x7    -> (sign extend) >> 1
//     // sra (sign) msb 0 // x8== 32'h0001_1000;
//     rom[8]  = 32'h40745433;
//     // slt x6, x10, x8   -> signed
//     // slt (Sign)  slt x6 , 
//     //x10(8000_0000) (-) < x8(0001_1000) (+)-> x6=1;
//     rom[9]  = 32'h00852333; 
//     // slt x6, x8, x10   -> signed
//      // slt (Sign) slt x6 , 
//      //x8(0001_1000) (+) < x10(8000_0000) (-) -> x6=0;
//     rom[10] = 32'h00A42333; 
//     // sltu x6, x10, x8  -> unsigned
//       // sltu (unsign)  slt x6 , 
//       //x10(msb==1) < x8(msb==0) -> x6=0;
//     rom[11] = 32'h00853333; 
//     // sltu x6, x8, x10  -> unsigned
//      // sltu (unsign) slt x6 , 
//      //x8(msb==0) < x10(msb==1) -> x6=1;
//     rom[12] = 32'h00A43333; 

//   end


// ---------------------------------------------------------------------------------------------------------------//
// ----------------------------------------------for_S-type-------------------------------------------------------//
// ---------------------------------------------------------------------------------------------------------------//

// initial begin
// // imm(7bit) , rs2(5bit)->x1 , rs1(5bit)->x2 , funct3(3bit) , imm(5bit) , op(7bit)
// // x1 = 32'h1111_1111 , x2 = 32'h2222_2222 , x3 =32'h3333_3333, x4=32'h4444_4444
// // x5 = 32'h2;
//     // ---------------- byte_off == 2'b00 ---------------- //
//         rom[0]  = 32'h0012A123; // sw x1, +2(x5)  [4] -> O
//         rom[1]  = 32'h00129323; // sh x1, +6(x5)  [8] -> O
//         rom[2]  = 32'h00128523; // sb x1, +10(x5) [12] -> O

//         // ---------------- byte_off == 2'b01 ---------------- //
//         rom[3]  = 32'h0022A1A3; // sw x2, +3(x5)  [5] -> X
//         rom[4]  = 32'h002293A3; // sh x2, +7(x5)  [9] -> X
//         rom[5]  = 32'h002285A3; // sb x2, +11(x5) [13] -> O

//         // ---------------- byte_off == 2'b10 ---------------- //
//         rom[6]  = 32'h0032A223; // sw x3, +4(x5)  [6] ->X
//         rom[7]  = 32'h00329423; // sh x3, +8(x5)  [10] ->O
//         rom[8]  = 32'h00328623; // sb x3, +12(x5) [14] ->O

//         // ---------------- byte_off == 2'b11 ---------------- //
//         rom[9]  = 32'h0042A2A3; // sw x4, +5(x5)  [7] -> X
//         rom[10] = 32'h004294A3; // sh x4, +9(x5)  [11] -> X
//         rom[11] = 32'h004286A3; // sb x4, +13(x5) [15] -> O
// end


// //---------------------------------------------------------------------------------------------------------------//
// //------------------------------------------------------for_IL_TYPE----------------------------------------------//
// //---------------------------------------------------------------------------------------------------------------//
    // initial begin
    //     //imm(12bit) rs1(5bit) funct3(3bit) rd(5bit) op(7bit)
    //     //data_mem[4]==32'h87654325
        
    //     // offset = 14 → imm = 14
    //     rom[0]  = 32'h00E12283; // lw  x5, 14(x2) -> O
    //     rom[1]  = 32'h00E11303; // lh  x6, 14(x2) -> O
    //     rom[2]  = 32'h00E10383; // lb  x7, 14(x2) -> O
    //     rom[3]  = 32'h00E15403; // lhu x8, 14(x2) -> O
    //     rom[4] = 32'h00E14483; // lbu x9, 14(x2) -> O

    //     // offset = 15 → imm = 15
    //     rom[5] = 32'h00F12283; // lw  x5, 15(x2) -> X
    //     rom[6] = 32'h00F11303; // lh  x6, 15(x2) -> X
    //     rom[7] = 32'h00F10383; // lb  x7, 15(x2) -> O
    //     rom[8] = 32'h00F15403; // lhu x8, 15(x2) -> X
    //     rom[9] = 32'h00F14483; // lbu x9, 15(x2) -> O

    //     // offset = 16 → imm = 16
    //     rom[10] = 32'h01012283; // lw  x5, 16(x2) -> X
    //     rom[11] = 32'h01011303; // lh  x6, 16(x2) -> O
    //     rom[12] = 32'h01010383; // lb  x7, 16(x2) -> O
    //     rom[13] = 32'h01015403; // lhu x8, 16(x2) -> O
    //     rom[14] = 32'h01014483; // lbu x9, 16(x2) -> O

    //     // offset = 17 → imm = 17
    //     rom[15] = 32'h01112283; // lw  x5, 17(x2) -> X
    //     rom[16] = 32'h01111303; // lh  x6, 17(x2) -> X
    //     rom[17] = 32'h01110383; // lb  x7, 17(x2) -> O
    //     rom[18] = 32'h01115403; // lhu x8, 17(x2) -> X
    //     rom[19] = 32'h01114483; // lbu x9, 17(x2) -> O



    // end
// //---------------------------------------------------------------------------------------------------------------//
// //------------------------------------------------for I_TYPE-----------------------------------------------------//
// //---------------------------------------------------------------------------------------------------------------//





    // initial begin
    //    //-------------------------------------I_TYPE--------------------------------------//
    //     //imm(12bit) rs1(5bit) funct3(3bit) rd(5bit) op(7bit)


    //     // I-type ALU & SHIFT (RV32I)
    //     rom[0] = 32'h00C5_0593;  // addi  x11, x10(10), 12                -> x11 <= 22
    //     rom[1] = 32'hFF45_0593;  // addi  x11, x10(10), -12               -> x11 <= -2
    //     rom[2] = 32'h00C6_A593;  // slti  x11, x13(13), 12                -> x11 <= 0 // signed compare
    //     rom[3] = 32'hFF46_A593;  // slti  x11, x13(13), -12               -> x11 <= 0
    //     rom[4] = 32'h00C6_B593;  // sltiu x11, x13(13), 0000_0000_1100    -> x11 <= 0 // unsigned compare
    //     rom[5] = 32'h080C_6B593; // sltiu x11, x13(13), 1000_0000_1100    -> x11 <= 1
    //     rom[6] = 32'h80C7_B593;  // sltiu x11, x15(8000_080C), 1000_0000_1100(0000_080C)    -> x11 <= 0
        

    //     rom[7] = 32'h0047_4593;  // xori  x11, x14(101), 4(100)           -> x11 <= 0b001
    //     rom[8] = 32'h0047_6593;  // ori   x11, x14(101), 4(100)           -> x11 <= 0b101
    //     rom[9] = 32'h0047_7593;  // andi  x11, x14(101), 4(100)           -> x11 <= 0b100

    //     // shift-immediates: imm[11:5]=funct7, imm[4:0]=shamt
    //     rom[10] = 32'h00C1_9593;  // slli  x11, x3(ffffffff), 12           -> 0xFFFF_FFFF << 12 = 0xFFFFF000
    //     rom[11] = 32'h00C1_D593;  // srli  x11, x3(ffffffff), 12           -> 0x000F_FFFF  // zero extended 
    //     rom[12] = 32'h40C1_D593;  // srai  x11, x3(ffffffff), 12           -> 0xFFFF_FFFF  // msb extended

    //     // try) inst_code[30]==1 
    //     // imm = 0100_0000_1100 (32'd1036) -> for add / for slt
    //     // imm = 1100_0000_1100  -> for slt
    //     // imm = 0100_0000_0100  -> for xor/and/or
    //     rom[13] = 32'h40C5_0593;  // addi  x11, x10(10), 0100_0000_1100     -> X11 <= 0x416
    //     rom[14] = 32'hC0C6_A593;  // slti  x11, x13(13), 1100_0000_1100(-)  -> X11 <= 0
    //     rom[15] = 32'h40C6_A593;  // slti  x11, x13(13), 0100_0000_1100(+)  -> X11 <= 1
    //     rom[16] = 32'hC0C6_B593;  // sltiu x11, x13(13), 1100_0000_1100(+)  -> X11 <= 1 
    //     rom[17] = 32'h40C6_B593;  // sltiu x11, x13(13), 0100_0000_1100(+)  -> X11 <= 1
    //     rom[18] = 32'h4047_4593;  // xori  x11, x14(101), 0100_0000_0100    -> X11 <= 0b0100_0000_0001
    //     rom[19] = 32'h4047_6593;  // ori   x11, x14(101), 0100_0000_0100    -> X11 <= 0b0100_0000_0101
    //     rom[20] = 32'h4047_7593;  // andi  x11, x14(101), 0100_0000_0100    -> X11 <= 0b0000_0000_0100
     
    // end


// //---------------------------------------------------------------------------------------------------------------//
// //------------------------------------------------for U_TYPE-----------------------------------------------------//
// //---------------------------------------------------------------------------------------------------------------//
//     initial begin       
//         // LUI rd imm20 // AUIP rd imm20
//           rom[0] = 32'hF00000B7; // LUI  x1,  20'hF0000   -> x1  <= 32'hF0000_000
//           rom[1] = 32'h10101137; // LUI  x2,  20'h10101   -> x2  <= 32'h10101_000
//           rom[2] = 32'hF0000197; // AUIPC x3, 20'hF0000   -> x3  <= 32'hF0000_000 + 32'd8
//           rom[3] = 32'h0000F217; // AUIPC x4, 20'h0000F   -> x4  <= 32'h0000F_000 + 32'd12
//           rom[4] = 32'h876542B7; // LUI  x5,  20'h87654   -> x5  <= 32'h87654_000
//           rom[5] = 32'h32128293; // ADDI x5, x5, 12'h321  -> x5  <= x5 + 0x321
//    end

// //---------------------------------------------------------------------------------------------------------------//
// //------------------------------------------------for JAL / JALR----------------------------------------------------//
// //---------------------------------------------------------------------------------------------------------------//
    // initial begin
    // // jal rd, offset        // rd = PC+4,   PC += offset
    // // jalr rd, rs1, imm12   // rd = PC+4,   PC = (rs1 + imm) & ~1

    // rom[0] = 32'h00C000EF; // pc=0   : jal  x1, +12   -> x1<=4,   PC<=12  (rom[3])             //[1]
    // rom[1] = 32'h00208133; // pc=4   : add  x2, x1, x2                                         //[4]
    // rom[2] = 32'h00C000EF; // pc=8   : jal  x1, +12   -> x1<=12,  PC<=20  (rom[5])             //[5]
    // rom[3] = 32'h00208133; // pc=12  : add  x2, x1, x2                                         //[2]
    // rom[4] = 32'h00008167; // pc=16  : jalr x2, x1, 0 -> x2<=20(0x14), PC<=x1(=4)  // return   //[3]
    // rom[5] = 32'hFEDFF0EF; // pc=20  : jal  x1, -20   -> 무한 루프 (PC=0)                       //[6] -> rom[0]
    // end



//---------------------------------------------sum=sum+a (a<11)-------------------------------------------------//
    // int a = 0;
    // int sum = 0;

    // while (a < 11) {      // 0~10 합: 55
    //     sum = adder(sum, a);
    //     a = a + 1;
    // }



//     x1 = ra (return address)
// x2 = sp (stack pointer)
// x5 = t0 (temporary)
// x8 = s0/fp (saved/frame pointer)
// x10 = a0, x11 = a1, x12 = a2, x13 = a3 (함수 인자/리턴)
// x18–x27 = s2–s11 (saved), x28–x31 = t3–t6 (temporaries)

    
    // initial begin
    //     // 0: sum=0;  1: a=0;
    //     rom[0]  = 32'h00000613; // addi x12, x0, 0      ; sum = 0
    //     rom[1]  = 32'h00000693; // addi x13, x0, 0      ; a   = 0

    //     // 2: t0 = (a < 11) ? 1:0
    //     rom[2]  = 32'h00b6a293; // slti x5, x13, 11

    //     // 3: if (t0 == 0) goto end(PC=40)
    //     rom[3]  = 32'h00028e63; // beq  x5, x0, +28     ; -> PC=40 (rom[10])
    //     // 4~6: a0=sum, a1=a, call adder
    //     rom[4]  = 32'h00060513; // addi x10, x12, 0     ; a0=sum
    //     rom[5]  = 32'h00068593; // addi x11, x13, 0     ; a1=a
    //     rom[6] = 32'h014000EF;  // jal x1, +20  (to rom[11])

    //     // 7: sum = return(a0);  8: a++
    //     rom[7]  = 32'h00050613; // addi x12, x10, 0     ; sum=a0
    //     rom[8]  = 32'h00168693; // addi x13, x13, 1     ; a=a+1

    //     // 9: goto loop(PC=8)
    //     rom[9] = 32'hFE5FF06F;  // jal x0, -28  (back to rom[2])

    //     // 10: end: 무한 대기
    //     rom[10] = 32'h0000006f; // jal  x0, 0           ; self-loop

    //     // 11~12: adder: a0 = a0 + a1; return
    //     rom[11] = 32'h00b50533; // add  x10, x10, x11   ; a0=a0+a1
    //     rom[12] = 32'h00008067; // jalr x0, x1, 0       ; ret
    // end






//-------------------------------------------------------------------------------------------------------------------------------//
    assign instr_code = rom[instr_rAddr[31:2]];

endmodule




//------------------------------------------b_type----------------------------------------------------------------//

// `timescale 1ns / 1ps

// module instr_mem (
//     input  logic [31:0] instr_rAddr,
//     output logic [31:0] instr_code
// );

//     logic [31:0] rom [0:63];

//     initial begin
//         for (int i = 0; i <64; i++) begin
//             rom[i] = 32'hffff_0000 + i;
//         end

//         rom[0] = 32'h004182B3; //32'b0000000_00100_00011_000_01010_0110011; // add x5, x3, x4
//         rom[1] = 32'h409403B3; //32'b0100000_01001_01000_000_01111_0110011; // sub x7, x8, x9

//         // B-type
//         // 32'b imm(7bit) _ rs2(5bit) _ rs1(5bit) _ funct3(3bit) _ imm(5bit) _ opcode(7'b1100011)
//         // rom[2] = 32'b0000000_00010_00010_000_10000_1100011;
//         rom[2] = 32'h00210863; // BEQ x2, x2, 16

//         // S-Type
//         // 32'b imm(7bit) _ rs2(5bit) _ rs1(5bit) _ funct3(3bit) _ imm(5bit) _ opcode(7'b0100011)
//         // rom[3] = 32'b0000000_00110_00100_010_00110_0100011;
//         rom[3] = 32'h00612323; // sb x6, 6(x2)
//         rom[4] = 32'h00811323; // sh x8, 6(x2)
//         rom[5] = 32'h00913223; // sw x9, 6(x2)
//         // 32'b0000000_00110_00100_010_00111_0100011
//         rom[6] = 32'h006103A3; // sb x6, 7(x2)

//         // IL-Type
//         // 32'b0000000_01100_01010_000_01100_0000011
//         rom[7] = 32'h00C12283; // lw x5, 12(x2)

//         // I-Type
//         // 32'b0000000_01000_01010_000_01100_0010011
//         rom[8] = 32'h00C30413; // addi x8, x6, 12
//     end
// assign instr_code = rom[instr_rAddr[31:2]];

// endmodule
